`timescale 1ns/1ps

/*
NANDy NAND gate CPU
*/

module nandy(
        input [7:0] ioain, iobin,
        output [7:0] ioaout, iobout,
        output brk
	);
endmodule